library verilog;
use verilog.vl_types.all;
entity ddr3 is
    generic(
        TCK_MIN         : integer := 1875;
        TJIT_PER        : integer := 90;
        TJIT_CC         : integer := 180;
        TERR_2PER       : integer := 132;
        TERR_3PER       : integer := 157;
        TERR_4PER       : integer := 175;
        TERR_5PER       : integer := 188;
        TERR_6PER       : integer := 200;
        TERR_7PER       : integer := 209;
        TERR_8PER       : integer := 217;
        TERR_9PER       : integer := 224;
        TERR_10PER      : integer := 231;
        TERR_11PER      : integer := 237;
        TERR_12PER      : integer := 242;
        TDS             : integer := 75;
        TDH             : integer := 100;
        TDQSQ           : integer := 150;
        TDQSS           : real    := 0.250000;
        TDSS            : real    := 0.200000;
        TDSH            : real    := 0.200000;
        TDQSCK          : integer := 300;
        TQSH            : real    := 0.380000;
        TQSL            : real    := 0.380000;
        TDIPW           : integer := 490;
        TIPW            : integer := 780;
        TIS             : integer := 275;
        TIH             : integer := 200;
        TRAS_MIN        : integer := 37500;
        TRC             : integer := 50625;
        TRCD            : integer := 13125;
        TRP             : integer := 13125;
        TXP             : integer := 7500;
        TCKE            : integer := 5625;
        TAON            : integer := 300;
        TWLS            : integer := 245;
        TWLH            : integer := 245;
        TWLO            : integer := 9000;
        TAA_MIN         : integer := 13125;
        CL_TIME         : integer := 13125;
        TRRD            : integer := 10000;
        TFAW            : integer := 50000;
        CL_MIN          : integer := 5;
        CL_MAX          : integer := 14;
        AL_MIN          : integer := 0;
        AL_MAX          : integer := 2;
        WR_MIN          : integer := 5;
        WR_MAX          : integer := 16;
        BL_MIN          : integer := 4;
        BL_MAX          : integer := 8;
        CWL_MIN         : integer := 5;
        CWL_MAX         : integer := 10;
        TCK_MAX         : integer := 3300;
        TCH_AVG_MIN     : real    := 0.470000;
        TCL_AVG_MIN     : real    := 0.470000;
        TCH_AVG_MAX     : real    := 0.530000;
        TCL_AVG_MAX     : real    := 0.530000;
        TCH_ABS_MIN     : real    := 0.430000;
        TCL_ABS_MIN     : real    := 0.430000;
        TCKE_TCK        : integer := 3;
        TAA_MAX         : integer := 20000;
        TQH             : real    := 0.380000;
        TRPRE           : real    := 0.900000;
        TRPST           : real    := 0.300000;
        TDQSH           : real    := 0.450000;
        TDQSL           : real    := 0.450000;
        TWPRE           : real    := 0.900000;
        TWPST           : real    := 0.300000;
        TZQCS           : integer := 64;
        TZQINIT         : integer := 512;
        TZQOPER         : integer := 256;
        TCCD            : integer := 4;
        TCCD_DG         : integer := 2;
        TRAS_MAX        : real    := 60000000000.000000;
        TWR             : integer := 15000;
        TMRD            : integer := 4;
        TMOD            : integer := 15000;
        TMOD_TCK        : integer := 12;
        TRRD_TCK        : integer := 4;
        TRRD_DG         : integer := 3000;
        TRRD_DG_TCK     : integer := 2;
        TRTP            : integer := 7500;
        TRTP_TCK        : integer := 4;
        TWTR            : integer := 7500;
        TWTR_DG         : integer := 3750;
        TWTR_TCK        : integer := 4;
        TWTR_DG_TCK     : integer := 2;
        TDLLK           : integer := 512;
        TRFC_MIN        : integer := 110000;
        TRFC_MAX        : integer := 70312500;
        TXP_TCK         : integer := 3;
        TXPDLL          : integer := 24000;
        TXPDLL_TCK      : integer := 10;
        TACTPDEN        : integer := 1;
        TPRPDEN         : integer := 1;
        TREFPDEN        : integer := 1;
        TCPDED          : integer := 1;
        TXPR            : integer := 120000;
        TXPR_TCK        : integer := 5;
        TXS             : integer := 120000;
        TXS_TCK         : integer := 5;
        TCKSRE          : integer := 10000;
        TCKSRE_TCK      : integer := 5;
        TCKSRX          : integer := 10000;
        TCKSRX_TCK      : integer := 5;
        TCKESR_TCK      : integer := 4;
        TAOF            : real    := 0.700000;
        TAONPD          : integer := 8500;
        TAOFPD          : integer := 8500;
        ODTH4           : integer := 4;
        ODTH8           : integer := 6;
        TADC            : real    := 0.700000;
        TWLMRD          : integer := 40;
        TWLDQSEN        : integer := 25;
        TWLOE           : integer := 2000;
        DM_BITS         : integer := 2;
        ADDR_BITS       : integer := 13;
        ROW_BITS        : integer := 13;
        COL_BITS        : integer := 10;
        DQ_BITS         : integer := 16;
        DQS_BITS        : integer := 2;
        BA_BITS         : integer := 3;
        MEM_BITS        : integer := 15;
        AP              : integer := 10;
        BC              : integer := 12;
        BL_BITS         : integer := 3;
        BO_BITS         : integer := 2;
        CS_BITS         : integer := 2;
        RANKS           : integer := 1;
        RZQ             : integer := 240;
        PRE_DEF_PAT     : integer := 170;
        STOP_ON_ERROR   : integer := 1;
        DEBUG           : integer := 0;
        BUS_DELAY       : integer := 0;
        RANDOM_OUT_DELAY: integer := 0;
        RANDOM_SEED     : integer := 711689044;
        RDQSEN_PRE      : integer := 2;
        RDQSEN_PST      : integer := 1;
        RDQS_PRE        : integer := 2;
        RDQS_PST        : integer := 1;
        RDQEN_PRE       : integer := 0;
        RDQEN_PST       : integer := 0;
        WDQS_PRE        : integer := 2;
        WDQS_PST        : integer := 1;
        check_strict_mrbits: integer := 1;
        check_strict_timing: integer := 1;
        feature_pasr    : integer := 1;
        feature_truebl4 : integer := 0;
        LOAD_MODE       : integer := 0;
        REFRESH         : integer := 1;
        PRECHARGE       : integer := 2;
        ACTIVATE        : integer := 3;
        WRITE           : integer := 4;
        READ            : integer := 5;
        ZQ              : integer := 6;
        NOP             : integer := 7;
        PWR_DOWN        : integer := 8;
        SELF_REF        : integer := 9;
        SAME_BANK       : integer := 0;
        DIFF_BANK       : integer := 1;
        DIFF_GROUP      : integer := 2
    );
    port(
        rst_n           : in     vl_logic;
        ck              : in     vl_logic;
        ck_n            : in     vl_logic;
        cke             : in     vl_logic;
        cs_n            : in     vl_logic;
        ras_n           : in     vl_logic;
        cas_n           : in     vl_logic;
        we_n            : in     vl_logic;
        dm_tdqs         : inout  vl_logic_vector;
        ba              : in     vl_logic_vector;
        addr            : in     vl_logic_vector;
        dq              : inout  vl_logic_vector;
        dqs             : inout  vl_logic_vector;
        dqs_n           : inout  vl_logic_vector;
        tdqs_n          : out    vl_logic_vector;
        odt             : in     vl_logic
    );
end ddr3;
